module vga_timing_top (
    input wire clk_100mhz,
    input wire clk_100mhz,
    output wire hsync,
    output wire vsync,
    output wire [7:0] rgb
);

pixel_clk_gen instance1 (

);

vga_timing_640x480 instance2 (

);