module vga_timing_640x480(
    input wire clk_pix,
    input wire clk_pix,
    output wire [9:0] hcount,
    output wire [9:0] hcount,
    output wire [9:0] hcount,
    output wire [9:0] hcount,
)